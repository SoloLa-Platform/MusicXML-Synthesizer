BZh91AY&SYS5�  �_�Px�ǟGװ?���@�N�Q��4�M� � 4h6�4H�	�S�4@  h �
�D�4ɽP  ���	DЩ�'�O)��&�f�F� �K�D
�X�C��Mi6�A�UɅ̣Ͷy,���l����>�L��g �U�^*�%��m�1������$�J���"��󲱡Zrn2��˧~Q)��pMcaBJ�T��N��J���-��(�n�!��>r����)Ď��c�E�)E�y�d����09H M�" ��~��|��A��e.h����mc{ }e"�\%��l
�b+�]IQ �:�)F�j�1\S��&�&����g�DE���*WX����$�h�D����%�M��`���K�"ª���n�B)��n/�sXp/q�Qz

��yB�A�dL�HV�L�'#��l�H�\T�����1T�P#T8:2�>�Ђ�B��]��BAL�0H